library ieee;
use ieee.std_logic_1164.all;
USE IEEE.numeric_std.ALL;

entity Instr_Memory is
  GENERIC (N:     NATURAL:= 32);  -- Width of inputs.
  port (address : in std_logic_vector(N-1 downto 0);			
		data    : out std_logic_vector(N-1 downto 0));
end Instr_Memory;

architecture behavioral of Instr_Memory is
signal addr : integer range 0 to 4*50760;  
 
begin
addr <= to_integer(unsigned(address));
   process(addr) 
	begin
      case addr is 
       when 4*0    => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*1    => data <= "10000110101000000000000000000001"; -- addi r21,r00,1
       when 4*2    => data <= "10000110110000000000000000000000"; -- addi r22,r00,0
       when 4*3    => data <= "10000100001000000000000000001010"; -- addi r01,r00,10
       when 4*4    => data <= "10000100010000000000000000001111"; -- addi r02,r00,15
       when 4*5    => data <= "10000100011000000000000000000101"; -- addi r03,r00,5
       when 4*6    => data <= "10000100100000000000000000000111"; -- addi r04,r00,7
       when 4*7    => data <= "10000100101000000000000000001100"; -- addi r05,r00,12
       when 4*8    => data <= "10000100110000000000000000010001"; -- addi r06,r00,17
       when 4*9    => data <= "10000100111000000000000000001101"; -- addi r07,r00,13
       when 4*10   => data <= "10000101000000000000000000000010"; -- addi r08,r00,2
       when 4*11   => data <= "00000000000000000000000000000000"; -- nop
       when 4*12   => data <= "00000000000000000000000000000000"; -- nop
       when 4*13   => data <= "00000000000000000000000000000000"; -- nop
       when 4*14   => data <= "00000000000000000000000000000000"; -- nop
       when 4*15   => data <= "00000000000000000000000000000000"; -- nop
       when 4*16   => data <= "11000000001000000000000000001011"; -- sb r01,r00,11
       when 4*17   => data <= "11000000010000000000000000001100"; -- sb r02,r00,12
       when 4*18   => data <= "11000000011000000000000000001101"; -- sb r03,r00,13
       when 4*19   => data <= "11000000100000000000000000001110"; -- sb r04,r00,14
       when 4*20   => data <= "11000000101000000000000000001111"; -- sb r05,r00,15
       when 4*21   => data <= "11000000110000000000000000010000"; -- sb r06,r00,16
       when 4*22   => data <= "11000000111000000000000000010001"; -- sb r07,r00,17
       when 4*23   => data <= "11000001000000000000000000010010"; -- sb r08,r00,18
       when 4*24   => data <= "00000000000000000000000000000000"; -- nop
       when 4*25   => data <= "00000000000000000000000000000000"; -- nop
       when 4*26   => data <= "00000000000000000000000000000000"; -- nop
       when 4*27   => data <= "00000000000000000000000000000000"; -- nop
       when 4*28   => data <= "00000000000000000000000000000000"; -- nop
       when 4*29   => data <= "10000101001000000000000000000110"; -- addi r09,r00,6
       when 4*30   => data <= "10000101010000000000000000000000"; -- addi r10,r00,0
       when 4*31   => data <= "10000101011000000000000000001000"; -- addi r11,r00,8
       when 4*32   => data <= "10000101100000000000000000000000"; -- addi r12,r00,0
       when 4*33   => data <= "00000000000000000000000000000000"; -- nop
       when 4*34   => data <= "00000000000000000000000000000000"; -- nop
       when 4*35   => data <= "00000000000000000000000000000000"; -- nop
       when 4*36   => data <= "00000000000000000000000000000000"; -- nop
       when 4*37   => data <= "00000000000000000000000000000000"; -- nop
       when 4*38   => data <= "10000000101010100000000000001011"; -- lb r05,r10,11
       when 4*39   => data <= "00000000000000000000000000000000"; -- nop
       when 4*40   => data <= "00000000000000000000000000000000"; -- nop
       when 4*41   => data <= "00000000000000000000000000000000"; -- nop
       when 4*42   => data <= "00000000000000000000000000000000"; -- nop
       when 4*43   => data <= "00000000000000000000000000000000"; -- nop
       when 4*44   => data <= "10000000110010100000000000001100"; -- lb r06,r10,12
       when 4*45   => data <= "00000000000000000000000000000000"; -- nop
       when 4*46   => data <= "00000000000000000000000000000000"; -- nop
       when 4*47   => data <= "00000000000000000000000000000000"; -- nop
       when 4*48   => data <= "00000000000000000000000000000000"; -- nop
       when 4*49   => data <= "00000000000000000000000000000000"; -- nop
       when 4*50   => data <= "10000100001001010000000000000000"; -- addi r01,r05,0
       when 4*51   => data <= "10000100010001100000000000000000"; -- addi r02,r06,0
       when 4*52   => data <= "00000000000000000000000000000000"; -- nop
       when 4*53   => data <= "00000000000000000000000000000000"; -- nop
       when 4*54   => data <= "00000000000000000000000000000000"; -- nop
       when 4*55   => data <= "00000000000000000000000000000000"; -- nop
       when 4*56   => data <= "00000000000000000000000000000000"; -- nop
       when 4*57   => data <= "00000000011000010001000000110100"; -- slt r03,r01,r02
       when 4*58   => data <= "00000000000000000000000000000000"; -- nop
       when 4*59   => data <= "00000000000000000000000000000000"; -- nop
       when 4*60   => data <= "00000000000000000000000000000000"; -- nop
       when 4*61   => data <= "00000000000000000000000000000000"; -- nop
       when 4*62   => data <= "00000000000000000000000000000000"; -- nop
       when 4*63   => data <= "00001000011000000000000001101011"; -- beq r03,r00,SWAP
       when 4*64   => data <= "00000000000000000000000000000000"; -- nop
       when 4*65   => data <= "00000000000000000000000000000000"; -- nop
       when 4*66   => data <= "00001001100010110000000111100110"; -- beq r12,r11,END
       when 4*67   => data <= "00000000000000000000000000000000"; -- nop
       when 4*68   => data <= "00000000000000000000000000000000"; -- nop
       when 4*69   => data <= "00000000000000000000000000000000"; -- nop
       when 4*70   => data <= "00000000000000000000000000000000"; -- nop
       when 4*71   => data <= "00000000000000000000000000000000"; -- nop
       when 4*72   => data <= "00001001010010010000000001001111"; -- beq r10,r09,INC2
       when 4*73   => data <= "00000000000000000000000000000000"; -- nop
       when 4*74   => data <= "00000000000000000000000000000000"; -- nop
       when 4*75   => data <= "00000000000000000000000000000000"; -- nop
       when 4*76   => data <= "00000100000000000000000001011110"; -- jmp INC1
       when 4*77   => data <= "00000000000000000000000000000000"; -- nop
       when 4*78   => data <= "00000000000000000000000000000000"; -- nop
       when 4*79   => data <= "00000000000000000000000000000000"; -- nop
       when 4*80   => data <= "00000000000000000000000000000000"; -- nop
       when 4*81   => data <= "00000000000000000000000000000000"; -- nop
       when 4*82   => data <= "10000101100011000000000000000001"; -- addi r12,r12,1
       when 4*83   => data <= "10000101010000000000000000000000"; -- addi r10,r00,0
       when 4*84   => data <= "10000110110000000000000000000000"; -- addi r22,r00,0
       when 4*85   => data <= "00000000000000000000000000000000"; -- nop
       when 4*86   => data <= "00000000000000000000000000000000"; -- nop
       when 4*87   => data <= "00000000000000000000000000000000"; -- nop
       when 4*88   => data <= "00000000000000000000000000000000"; -- nop
       when 4*89   => data <= "00000000000000000000000000000000"; -- nop
       when 4*90   => data <= "00000100000000000000000001111100"; -- jmp OUTPUT
       when 4*91   => data <= "00000000000000000000000000000000"; -- nop
       when 4*92   => data <= "00000000000000000000000000000000"; -- nop
       when 4*93   => data <= "00000000000000000000000000000000"; -- nop
       when 4*94   => data <= "00000000000000000000000000000000"; -- nop
       when 4*95   => data <= "00000000000000000000000000000000"; -- nop
       when 4*96   => data <= "00000000000000000000000000000000"; -- nop
       when 4*97   => data <= "00000000000000000000000000000000"; -- nop
       when 4*98   => data <= "10000101010010100000000000000001"; -- addi r10,r10,1
       when 4*99   => data <= "00000000000000000000000000000000"; -- nop
       when 4*100   => data <= "00000000000000000000000000000000"; -- nop
       when 4*101   => data <= "00000000000000000000000000000000"; -- nop
       when 4*102   => data <= "00000000000000000000000000000000"; -- nop
       when 4*103   => data <= "00000000000000000000000000000000"; -- nop
       when 4*104   => data <= "00000100000000000000000000100001"; -- jmp LOOP
       when 4*105   => data <= "00000000000000000000000000000000"; -- nop
       when 4*106   => data <= "00000000000000000000000000000000"; -- nop
       when 4*107   => data <= "00000000000000000000000000000000"; -- nop
       when 4*108   => data <= "00000000000000000000000000000000"; -- nop
       when 4*109   => data <= "00000000000000000000000000000000"; -- nop
       when 4*110   => data <= "00000000000000000000000000000000"; -- nop
       when 4*111   => data <= "00000000000000000000000000000000"; -- nop
       when 4*112   => data <= "11000000010010100000000000001011"; -- sb r02,r10,11
       when 4*113   => data <= "00000000000000000000000000000000"; -- nop
       when 4*114   => data <= "00000000000000000000000000000000"; -- nop
       when 4*115   => data <= "11000000001010100000000000001100"; -- sb r01,r10,12
       when 4*116   => data <= "00000000000000000000000000000000"; -- nop
       when 4*117   => data <= "00000000000000000000000000000000"; -- nop
       when 4*118   => data <= "00000000000000000000000000000000"; -- nop
       when 4*119   => data <= "00000000000000000000000000000000"; -- nop
       when 4*120   => data <= "00000000000000000000000000000000"; -- nop
       when 4*121   => data <= "00000100000000000000000001000010"; -- jmp SWAPPED
       when 4*122   => data <= "00000000000000000000000000000000"; -- nop
       when 4*123   => data <= "00000000000000000000000000000000"; -- nop
       when 4*124   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*125   => data <= "00000000000000000000000000000000"; -- nop
       when 4*126   => data <= "00000000000000000000000000000000"; -- nop
       when 4*127   => data <= "00000000000000000000000000000000"; -- nop
       when 4*128   => data <= "00000000000000000000000000000000"; -- nop
       when 4*129   => data <= "00000000000000000000000000000000"; -- nop
       when 4*130   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*131   => data <= "00000000000000000000000000000000"; -- nop
       when 4*132   => data <= "00000000000000000000000000000000"; -- nop
       when 4*133   => data <= "00000000000000000000000000000000"; -- nop
       when 4*134   => data <= "00000000000000000000000000000000"; -- nop
       when 4*135   => data <= "00000000000000000000000000000000"; -- nop
       when 4*136   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*137   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*138   => data <= "00000100000000000000000100011110"; -- jmp LOOP1
       when 4*139   => data <= "00000000000000000000000000000000"; -- nop
       when 4*140   => data <= "00000000000000000000000000000000"; -- nop
       when 4*141   => data <= "00000000000000000000000000000000"; -- nop
       when 4*142   => data <= "00000000000000000000000000000000"; -- nop
       when 4*143   => data <= "00000000000000000000000000000000"; -- nop
       when 4*144   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*145   => data <= "00000000000000000000000000000000"; -- nop
       when 4*146   => data <= "00000000000000000000000000000000"; -- nop
       when 4*147   => data <= "00000000000000000000000000000000"; -- nop
       when 4*148   => data <= "00000000000000000000000000000000"; -- nop
       when 4*149   => data <= "00000000000000000000000000000000"; -- nop
       when 4*150   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*151   => data <= "00000000000000000000000000000000"; -- nop
       when 4*152   => data <= "00000000000000000000000000000000"; -- nop
       when 4*153   => data <= "00000000000000000000000000000000"; -- nop
       when 4*154   => data <= "00000000000000000000000000000000"; -- nop
       when 4*155   => data <= "00000000000000000000000000000000"; -- nop
       when 4*156   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*157   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*158   => data <= "00000100000000000000000100110111"; -- jmp LOOP2
       when 4*159   => data <= "00000000000000000000000000000000"; -- nop
       when 4*160   => data <= "00000000000000000000000000000000"; -- nop
       when 4*161   => data <= "00000000000000000000000000000000"; -- nop
       when 4*162   => data <= "00000000000000000000000000000000"; -- nop
       when 4*163   => data <= "00000000000000000000000000000000"; -- nop
       when 4*164   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*165   => data <= "00000000000000000000000000000000"; -- nop
       when 4*166   => data <= "00000000000000000000000000000000"; -- nop
       when 4*167   => data <= "00000000000000000000000000000000"; -- nop
       when 4*168   => data <= "00000000000000000000000000000000"; -- nop
       when 4*169   => data <= "00000000000000000000000000000000"; -- nop
       when 4*170   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*171   => data <= "00000000000000000000000000000000"; -- nop
       when 4*172   => data <= "00000000000000000000000000000000"; -- nop
       when 4*173   => data <= "00000000000000000000000000000000"; -- nop
       when 4*174   => data <= "00000000000000000000000000000000"; -- nop
       when 4*175   => data <= "00000000000000000000000000000000"; -- nop
       when 4*176   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*177   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*178   => data <= "00000100000000000000000101010000"; -- jmp LOOP3
       when 4*179   => data <= "00000000000000000000000000000000"; -- nop
       when 4*180   => data <= "00000000000000000000000000000000"; -- nop
       when 4*181   => data <= "00000000000000000000000000000000"; -- nop
       when 4*182   => data <= "00000000000000000000000000000000"; -- nop
       when 4*183   => data <= "00000000000000000000000000000000"; -- nop
       when 4*184   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*185   => data <= "00000000000000000000000000000000"; -- nop
       when 4*186   => data <= "00000000000000000000000000000000"; -- nop
       when 4*187   => data <= "00000000000000000000000000000000"; -- nop
       when 4*188   => data <= "00000000000000000000000000000000"; -- nop
       when 4*189   => data <= "00000000000000000000000000000000"; -- nop
       when 4*190   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*191   => data <= "00000000000000000000000000000000"; -- nop
       when 4*192   => data <= "00000000000000000000000000000000"; -- nop
       when 4*193   => data <= "00000000000000000000000000000000"; -- nop
       when 4*194   => data <= "00000000000000000000000000000000"; -- nop
       when 4*195   => data <= "00000000000000000000000000000000"; -- nop
       when 4*196   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*197   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*198   => data <= "00000100000000000000000101101001"; -- jmp LOOP4
       when 4*199   => data <= "00000000000000000000000000000000"; -- nop
       when 4*200   => data <= "00000000000000000000000000000000"; -- nop
       when 4*201   => data <= "00000000000000000000000000000000"; -- nop
       when 4*202   => data <= "00000000000000000000000000000000"; -- nop
       when 4*203   => data <= "00000000000000000000000000000000"; -- nop
       when 4*204   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*205   => data <= "00000000000000000000000000000000"; -- nop
       when 4*206   => data <= "00000000000000000000000000000000"; -- nop
       when 4*207   => data <= "00000000000000000000000000000000"; -- nop
       when 4*208   => data <= "00000000000000000000000000000000"; -- nop
       when 4*209   => data <= "00000000000000000000000000000000"; -- nop
       when 4*210   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*211   => data <= "00000000000000000000000000000000"; -- nop
       when 4*212   => data <= "00000000000000000000000000000000"; -- nop
       when 4*213   => data <= "00000000000000000000000000000000"; -- nop
       when 4*214   => data <= "00000000000000000000000000000000"; -- nop
       when 4*215   => data <= "00000000000000000000000000000000"; -- nop
       when 4*216   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*217   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*218   => data <= "00000100000000000000000110000010"; -- jmp LOOP5
       when 4*219   => data <= "00000000000000000000000000000000"; -- nop
       when 4*220   => data <= "00000000000000000000000000000000"; -- nop
       when 4*221   => data <= "00000000000000000000000000000000"; -- nop
       when 4*222   => data <= "00000000000000000000000000000000"; -- nop
       when 4*223   => data <= "00000000000000000000000000000000"; -- nop
       when 4*224   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*225   => data <= "00000000000000000000000000000000"; -- nop
       when 4*226   => data <= "00000000000000000000000000000000"; -- nop
       when 4*227   => data <= "00000000000000000000000000000000"; -- nop
       when 4*228   => data <= "00000000000000000000000000000000"; -- nop
       when 4*229   => data <= "00000000000000000000000000000000"; -- nop
       when 4*230   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*231   => data <= "00000000000000000000000000000000"; -- nop
       when 4*232   => data <= "00000000000000000000000000000000"; -- nop
       when 4*233   => data <= "00000000000000000000000000000000"; -- nop
       when 4*234   => data <= "00000000000000000000000000000000"; -- nop
       when 4*235   => data <= "00000000000000000000000000000000"; -- nop
       when 4*236   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*237   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*238   => data <= "00000100000000000000000110011011"; -- jmp LOOP6
       when 4*239   => data <= "00000000000000000000000000000000"; -- nop
       when 4*240   => data <= "00000000000000000000000000000000"; -- nop
       when 4*241   => data <= "00000000000000000000000000000000"; -- nop
       when 4*242   => data <= "00000000000000000000000000000000"; -- nop
       when 4*243   => data <= "00000000000000000000000000000000"; -- nop
       when 4*244   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*245   => data <= "00000000000000000000000000000000"; -- nop
       when 4*246   => data <= "00000000000000000000000000000000"; -- nop
       when 4*247   => data <= "00000000000000000000000000000000"; -- nop
       when 4*248   => data <= "00000000000000000000000000000000"; -- nop
       when 4*249   => data <= "00000000000000000000000000000000"; -- nop
       when 4*250   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*251   => data <= "00000000000000000000000000000000"; -- nop
       when 4*252   => data <= "00000000000000000000000000000000"; -- nop
       when 4*253   => data <= "00000000000000000000000000000000"; -- nop
       when 4*254   => data <= "00000000000000000000000000000000"; -- nop
       when 4*255   => data <= "00000000000000000000000000000000"; -- nop
       when 4*256   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*257   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*258   => data <= "00000100000000000000000110110100"; -- jmp LOOP7
       when 4*259   => data <= "00000000000000000000000000000000"; -- nop
       when 4*260   => data <= "00000000000000000000000000000000"; -- nop
       when 4*261   => data <= "00000000000000000000000000000000"; -- nop
       when 4*262   => data <= "00000000000000000000000000000000"; -- nop
       when 4*263   => data <= "00000000000000000000000000000000"; -- nop
       when 4*264   => data <= "10000110110101100000000000000001"; -- addi r22,r22,1
       when 4*265   => data <= "00000000000000000000000000000000"; -- nop
       when 4*266   => data <= "00000000000000000000000000000000"; -- nop
       when 4*267   => data <= "00000000000000000000000000000000"; -- nop
       when 4*268   => data <= "00000000000000000000000000000000"; -- nop
       when 4*269   => data <= "00000000000000000000000000000000"; -- nop
       when 4*270   => data <= "10000011110101100000000000001010"; -- lb r30,r22,10
       when 4*271   => data <= "00000000000000000000000000000000"; -- nop
       when 4*272   => data <= "00000000000000000000000000000000"; -- nop
       when 4*273   => data <= "00000000000000000000000000000000"; -- nop
       when 4*274   => data <= "00000000000000000000000000000000"; -- nop
       when 4*275   => data <= "00000000000000000000000000000000"; -- nop
       when 4*276   => data <= "10000110100000000000000000000010"; -- addi r20,r00,2
       when 4*277   => data <= "11000011110000000000000000000000"; -- sb r30,r00,0
       when 4*278   => data <= "00000100000000000000000111001101"; -- jmp LOOP8
       when 4*279   => data <= "00000000000000000000000000000000"; -- nop
       when 4*280   => data <= "00000000000000000000000000000000"; -- nop
       when 4*281   => data <= "00000000000000000000000000000000"; -- nop
       when 4*282   => data <= "00000000000000000000000000000000"; -- nop
       when 4*283   => data <= "00000000000000000000000000000000"; -- nop
       when 4*284   => data <= "00000000000000000000000000000000"; -- nop
       when 4*285   => data <= "00000000000000000000000000000000"; -- nop
       when 4*286   => data <= "00001010100000000000000010010000"; -- beq r20,r00,O2
       when 4*287   => data <= "00000000000000000000000000000000"; -- nop
       when 4*288   => data <= "00000000000000000000000000000000"; -- nop
       when 4*289   => data <= "00000000000000000000000000000000"; -- nop
       when 4*290   => data <= "00000000000000000000000000000000"; -- nop
       when 4*291   => data <= "00000000000000000000000000000000"; -- nop
       when 4*292   => data <= "00000000000000000000000000000000"; -- nop
       when 4*293   => data <= "00000000000000000000000000000000"; -- nop
       when 4*294   => data <= "00000000000000000000000000000000"; -- nop
       when 4*295   => data <= "00000000000000000000000000000000"; -- nop
       when 4*296   => data <= "00000000000000000000000000000000"; -- nop
       when 4*297   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*298   => data <= "00000000000000000000000000000000"; -- nop
       when 4*299   => data <= "00000000000000000000000000000000"; -- nop
       when 4*300   => data <= "00000000000000000000000000000000"; -- nop
       when 4*301   => data <= "00000000000000000000000000000000"; -- nop
       when 4*302   => data <= "00000000000000000000000000000000"; -- nop
       when 4*303   => data <= "00000000000000000000000000000000"; -- nop
       when 4*304   => data <= "00000000000000000000000000000000"; -- nop
       when 4*305   => data <= "00000000000000000000000000000000"; -- nop
       when 4*306   => data <= "00000000000000000000000000000000"; -- nop
       when 4*307   => data <= "00000000000000000000000000000000"; -- nop
       when 4*308   => data <= "00000100000000000000000100011110"; -- jmp LOOP1
       when 4*309   => data <= "00000000000000000000000000000000"; -- nop
       when 4*310   => data <= "00000000000000000000000000000000"; -- nop
       when 4*311   => data <= "00001010100000000000000010100100"; -- beq r20,r00,O3
       when 4*312   => data <= "00000000000000000000000000000000"; -- nop
       when 4*313   => data <= "00000000000000000000000000000000"; -- nop
       when 4*314   => data <= "00000000000000000000000000000000"; -- nop
       when 4*315   => data <= "00000000000000000000000000000000"; -- nop
       when 4*316   => data <= "00000000000000000000000000000000"; -- nop
       when 4*317   => data <= "00000000000000000000000000000000"; -- nop
       when 4*318   => data <= "00000000000000000000000000000000"; -- nop
       when 4*319   => data <= "00000000000000000000000000000000"; -- nop
       when 4*320   => data <= "00000000000000000000000000000000"; -- nop
       when 4*321   => data <= "00000000000000000000000000000000"; -- nop
       when 4*322   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*323   => data <= "00000000000000000000000000000000"; -- nop
       when 4*324   => data <= "00000000000000000000000000000000"; -- nop
       when 4*325   => data <= "00000000000000000000000000000000"; -- nop
       when 4*326   => data <= "00000000000000000000000000000000"; -- nop
       when 4*327   => data <= "00000000000000000000000000000000"; -- nop
       when 4*328   => data <= "00000000000000000000000000000000"; -- nop
       when 4*329   => data <= "00000000000000000000000000000000"; -- nop
       when 4*330   => data <= "00000000000000000000000000000000"; -- nop
       when 4*331   => data <= "00000000000000000000000000000000"; -- nop
       when 4*332   => data <= "00000000000000000000000000000000"; -- nop
       when 4*333   => data <= "00000100000000000000000100110111"; -- jmp LOOP2
       when 4*334   => data <= "00000000000000000000000000000000"; -- nop
       when 4*335   => data <= "00000000000000000000000000000000"; -- nop
       when 4*336   => data <= "00001010100000000000000010111000"; -- beq r20,r00,O4
       when 4*337   => data <= "00000000000000000000000000000000"; -- nop
       when 4*338   => data <= "00000000000000000000000000000000"; -- nop
       when 4*339   => data <= "00000000000000000000000000000000"; -- nop
       when 4*340   => data <= "00000000000000000000000000000000"; -- nop
       when 4*341   => data <= "00000000000000000000000000000000"; -- nop
       when 4*342   => data <= "00000000000000000000000000000000"; -- nop
       when 4*343   => data <= "00000000000000000000000000000000"; -- nop
       when 4*344   => data <= "00000000000000000000000000000000"; -- nop
       when 4*345   => data <= "00000000000000000000000000000000"; -- nop
       when 4*346   => data <= "00000000000000000000000000000000"; -- nop
       when 4*347   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*348   => data <= "00000000000000000000000000000000"; -- nop
       when 4*349   => data <= "00000000000000000000000000000000"; -- nop
       when 4*350   => data <= "00000000000000000000000000000000"; -- nop
       when 4*351   => data <= "00000000000000000000000000000000"; -- nop
       when 4*352   => data <= "00000000000000000000000000000000"; -- nop
       when 4*353   => data <= "00000000000000000000000000000000"; -- nop
       when 4*354   => data <= "00000000000000000000000000000000"; -- nop
       when 4*355   => data <= "00000000000000000000000000000000"; -- nop
       when 4*356   => data <= "00000000000000000000000000000000"; -- nop
       when 4*357   => data <= "00000000000000000000000000000000"; -- nop
       when 4*358   => data <= "00000100000000000000000101010000"; -- jmp LOOP3
       when 4*359   => data <= "00000000000000000000000000000000"; -- nop
       when 4*360   => data <= "00000000000000000000000000000000"; -- nop
       when 4*361   => data <= "00001010100000000000000011001100"; -- beq r20,r00,O5
       when 4*362   => data <= "00000000000000000000000000000000"; -- nop
       when 4*363   => data <= "00000000000000000000000000000000"; -- nop
       when 4*364   => data <= "00000000000000000000000000000000"; -- nop
       when 4*365   => data <= "00000000000000000000000000000000"; -- nop
       when 4*366   => data <= "00000000000000000000000000000000"; -- nop
       when 4*367   => data <= "00000000000000000000000000000000"; -- nop
       when 4*368   => data <= "00000000000000000000000000000000"; -- nop
       when 4*369   => data <= "00000000000000000000000000000000"; -- nop
       when 4*370   => data <= "00000000000000000000000000000000"; -- nop
       when 4*371   => data <= "00000000000000000000000000000000"; -- nop
       when 4*372   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*373   => data <= "00000000000000000000000000000000"; -- nop
       when 4*374   => data <= "00000000000000000000000000000000"; -- nop
       when 4*375   => data <= "00000000000000000000000000000000"; -- nop
       when 4*376   => data <= "00000000000000000000000000000000"; -- nop
       when 4*377   => data <= "00000000000000000000000000000000"; -- nop
       when 4*378   => data <= "00000000000000000000000000000000"; -- nop
       when 4*379   => data <= "00000000000000000000000000000000"; -- nop
       when 4*380   => data <= "00000000000000000000000000000000"; -- nop
       when 4*381   => data <= "00000000000000000000000000000000"; -- nop
       when 4*382   => data <= "00000000000000000000000000000000"; -- nop
       when 4*383   => data <= "00000100000000000000000101101001"; -- jmp LOOP4
       when 4*384   => data <= "00000000000000000000000000000000"; -- nop
       when 4*385   => data <= "00000000000000000000000000000000"; -- nop
       when 4*386   => data <= "00001010100000000000000011100000"; -- beq r20,r00,O6
       when 4*387   => data <= "00000000000000000000000000000000"; -- nop
       when 4*388   => data <= "00000000000000000000000000000000"; -- nop
       when 4*389   => data <= "00000000000000000000000000000000"; -- nop
       when 4*390   => data <= "00000000000000000000000000000000"; -- nop
       when 4*391   => data <= "00000000000000000000000000000000"; -- nop
       when 4*392   => data <= "00000000000000000000000000000000"; -- nop
       when 4*393   => data <= "00000000000000000000000000000000"; -- nop
       when 4*394   => data <= "00000000000000000000000000000000"; -- nop
       when 4*395   => data <= "00000000000000000000000000000000"; -- nop
       when 4*396   => data <= "00000000000000000000000000000000"; -- nop
       when 4*397   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*398   => data <= "00000000000000000000000000000000"; -- nop
       when 4*399   => data <= "00000000000000000000000000000000"; -- nop
       when 4*400   => data <= "00000000000000000000000000000000"; -- nop
       when 4*401   => data <= "00000000000000000000000000000000"; -- nop
       when 4*402   => data <= "00000000000000000000000000000000"; -- nop
       when 4*403   => data <= "00000000000000000000000000000000"; -- nop
       when 4*404   => data <= "00000000000000000000000000000000"; -- nop
       when 4*405   => data <= "00000000000000000000000000000000"; -- nop
       when 4*406   => data <= "00000000000000000000000000000000"; -- nop
       when 4*407   => data <= "00000000000000000000000000000000"; -- nop
       when 4*408   => data <= "00000100000000000000000110000010"; -- jmp LOOP5
       when 4*409   => data <= "00000000000000000000000000000000"; -- nop
       when 4*410   => data <= "00000000000000000000000000000000"; -- nop
       when 4*411   => data <= "00001010100000000000000011110100"; -- beq r20,r00,O7
       when 4*412   => data <= "00000000000000000000000000000000"; -- nop
       when 4*413   => data <= "00000000000000000000000000000000"; -- nop
       when 4*414   => data <= "00000000000000000000000000000000"; -- nop
       when 4*415   => data <= "00000000000000000000000000000000"; -- nop
       when 4*416   => data <= "00000000000000000000000000000000"; -- nop
       when 4*417   => data <= "00000000000000000000000000000000"; -- nop
       when 4*418   => data <= "00000000000000000000000000000000"; -- nop
       when 4*419   => data <= "00000000000000000000000000000000"; -- nop
       when 4*420   => data <= "00000000000000000000000000000000"; -- nop
       when 4*421   => data <= "00000000000000000000000000000000"; -- nop
       when 4*422   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*423   => data <= "00000000000000000000000000000000"; -- nop
       when 4*424   => data <= "00000000000000000000000000000000"; -- nop
       when 4*425   => data <= "00000000000000000000000000000000"; -- nop
       when 4*426   => data <= "00000000000000000000000000000000"; -- nop
       when 4*427   => data <= "00000000000000000000000000000000"; -- nop
       when 4*428   => data <= "00000000000000000000000000000000"; -- nop
       when 4*429   => data <= "00000000000000000000000000000000"; -- nop
       when 4*430   => data <= "00000000000000000000000000000000"; -- nop
       when 4*431   => data <= "00000000000000000000000000000000"; -- nop
       when 4*432   => data <= "00000000000000000000000000000000"; -- nop
       when 4*433   => data <= "00000100000000000000000110011011"; -- jmp LOOP6
       when 4*434   => data <= "00000000000000000000000000000000"; -- nop
       when 4*435   => data <= "00000000000000000000000000000000"; -- nop
       when 4*436   => data <= "00001010100000000000000100001000"; -- beq r20,r00,O8
       when 4*437   => data <= "00000000000000000000000000000000"; -- nop
       when 4*438   => data <= "00000000000000000000000000000000"; -- nop
       when 4*439   => data <= "00000000000000000000000000000000"; -- nop
       when 4*440   => data <= "00000000000000000000000000000000"; -- nop
       when 4*441   => data <= "00000000000000000000000000000000"; -- nop
       when 4*442   => data <= "00000000000000000000000000000000"; -- nop
       when 4*443   => data <= "00000000000000000000000000000000"; -- nop
       when 4*444   => data <= "00000000000000000000000000000000"; -- nop
       when 4*445   => data <= "00000000000000000000000000000000"; -- nop
       when 4*446   => data <= "00000000000000000000000000000000"; -- nop
       when 4*447   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*448   => data <= "00000000000000000000000000000000"; -- nop
       when 4*449   => data <= "00000000000000000000000000000000"; -- nop
       when 4*450   => data <= "00000000000000000000000000000000"; -- nop
       when 4*451   => data <= "00000000000000000000000000000000"; -- nop
       when 4*452   => data <= "00000000000000000000000000000000"; -- nop
       when 4*453   => data <= "00000000000000000000000000000000"; -- nop
       when 4*454   => data <= "00000000000000000000000000000000"; -- nop
       when 4*455   => data <= "00000000000000000000000000000000"; -- nop
       when 4*456   => data <= "00000000000000000000000000000000"; -- nop
       when 4*457   => data <= "00000000000000000000000000000000"; -- nop
       when 4*458   => data <= "00000100000000000000000110110100"; -- jmp LOOP7
       when 4*459   => data <= "00000000000000000000000000000000"; -- nop
       when 4*460   => data <= "00000000000000000000000000000000"; -- nop
       when 4*461   => data <= "00001010100000000000000000100001"; -- beq r20,r00,LOOP
       when 4*462   => data <= "00000000000000000000000000000000"; -- nop
       when 4*463   => data <= "00000000000000000000000000000000"; -- nop
       when 4*464   => data <= "00000000000000000000000000000000"; -- nop
       when 4*465   => data <= "00000000000000000000000000000000"; -- nop
       when 4*466   => data <= "00000000000000000000000000000000"; -- nop
       when 4*467   => data <= "00000000000000000000000000000000"; -- nop
       when 4*468   => data <= "00000000000000000000000000000000"; -- nop
       when 4*469   => data <= "00000000000000000000000000000000"; -- nop
       when 4*470   => data <= "00000000000000000000000000000000"; -- nop
       when 4*471   => data <= "00000000000000000000000000000000"; -- nop
       when 4*472   => data <= "00000010100101001010100000100010"; -- sub r20,r20,r21
       when 4*473   => data <= "00000000000000000000000000000000"; -- nop
       when 4*474   => data <= "00000000000000000000000000000000"; -- nop
       when 4*475   => data <= "00000000000000000000000000000000"; -- nop
       when 4*476   => data <= "00000000000000000000000000000000"; -- nop
       when 4*477   => data <= "00000000000000000000000000000000"; -- nop
       when 4*478   => data <= "00000000000000000000000000000000"; -- nop
       when 4*479   => data <= "00000000000000000000000000000000"; -- nop
       when 4*480   => data <= "00000000000000000000000000000000"; -- nop
       when 4*481   => data <= "00000000000000000000000000000000"; -- nop
       when 4*482   => data <= "00000000000000000000000000000000"; -- nop
       when 4*483   => data <= "00000100000000000000000111001101"; -- jmp LOOP8
       when 4*484   => data <= "00000000000000000000000000000000"; -- nop
       when 4*485   => data <= "00000000000000000000000000000000"; -- nop
       when 4*486   => data <= "00000000000000000000000000000000"; -- nop
       when 4*487   => data <= "00000000000000000000000000000000"; -- nop
       when 4*488   => data <= "00000000000000000000000000000000"; -- nop
	    when others => data <= "00000000000000000000000000000000"; 
       end case;
	end process;
end behavioral;
