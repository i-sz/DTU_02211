library ieee;
use ieee.std_logic_1164.all;
USE IEEE.numeric_std.ALL;

entity Instr_Memory is
  GENERIC (N:     NATURAL:= 32);  -- Width of inputs.
  port (address : in std_logic_vector(N-1 downto 0);			
		data    : out std_logic_vector(N-1 downto 0));
end Instr_Memory;

architecture behavioral of Instr_Memory is
signal addr : integer range 0 to 4*50760;  
 
begin
addr <= to_integer(unsigned(address));
   process(addr) 
	begin
      case addr is 
       when 4*0    => data <= "00000000000000000000000000000000"; -- nop
       when 4*1    => data <= "10000100001000010000000000001010"; -- addi r01,r01,10
       when 4*2    => data <= "00000000000000000000000000000000"; -- nop
       when 4*3    => data <= "10000100010000000000000000000000"; -- addi r02,r00,0
       when 4*4    => data <= "00000000000000000000000000000000"; -- nop
       when 4*5    => data <= "00000000000000000000000000000000"; -- nop
       when 4*6    => data <= "00000000000000000000000000000000"; -- nop
       when 4*7    => data <= "00000000000000000000000000000000"; -- nop
       when 4*8    => data <= "00000000000000000000000000000000"; -- nop
       when 4*9    => data <= "00001000001000100000000000010110"; -- beq r01,r02,LOOP2IN
       when 4*10   => data <= "00000000000000000000000000000000"; -- nop
       when 4*11   => data <= "00000000000000000000000000000000"; -- nop
       when 4*12   => data <= "00000000000000000000000000000000"; -- nop
       when 4*13   => data <= "00000000000000000000000000000000"; -- nop
       when 4*14   => data <= "00000000000000000000000000000000"; -- nop
       when 4*15   => data <= "11000000010000100000000000000000"; -- sb r02,r02,0
       when 4*16   => data <= "10000100010000100000000000000001"; -- addi r02,r02,1
       when 4*17   => data <= "00000000000000000000000000000000"; -- nop
       when 4*18   => data <= "00000100000000000000000000001001"; -- jmp LOOP
       when 4*19   => data <= "00000000000000000000000000000000"; -- nop
       when 4*20   => data <= "00000000000000000000000000000000"; -- nop
       when 4*21   => data <= "00000000000000000000000000000000"; -- nop
       when 4*22   => data <= "10000100011000100000000000000000"; -- addi r03,r02,0
       when 4*23   => data <= "10000100010000000000000000000000"; -- addi r02,r00,0
       when 4*24   => data <= "00000000000000000000000000000000"; -- nop
       when 4*25   => data <= "00000000000000000000000000000000"; -- nop
       when 4*26   => data <= "00000000000000000000000000000000"; -- nop
       when 4*27   => data <= "00000000000000000000000000000000"; -- nop
       when 4*28   => data <= "00000000000000000000000000000000"; -- nop
       when 4*29   => data <= "00001000010000110000000000101011"; -- beq r02,r03,END
       when 4*30   => data <= "00000000000000000000000000000000"; -- nop
       when 4*31   => data <= "00000000000000000000000000000000"; -- nop
       when 4*32   => data <= "00000000000000000000000000000000"; -- nop
       when 4*33   => data <= "00000000000000000000000000000000"; -- nop
       when 4*34   => data <= "00000000000000000000000000000000"; -- nop
       when 4*35   => data <= "10000000100000100000000000000000"; -- lb r04,r02,0
       when 4*36   => data <= "10000100010000100000000000000001"; -- addi r02,r02,1
       when 4*37   => data <= "00000000000000000000000000000000"; -- nop
       when 4*38   => data <= "00000000000000000000000000000000"; -- nop
       when 4*39   => data <= "00000000000000000000000000000000"; -- nop
       when 4*40   => data <= "00000100000000000000000000011101"; -- jmp LOOP2
       when 4*41   => data <= "00000000000000000000000000000000"; -- nop
       when 4*42   => data <= "00000000000000000000000000000000"; -- nop
       when 4*43   => data <= "00000000000000000000000000000000"; -- nop
       when 4*44   => data <= "00000000000000000000000000000000"; -- nop
	    when others => data <= "00000000000000000000000000000000"; 
       end case;
	end process;
end behavioral;
