library ieee;
use ieee.std_logic_1164.all;
USE IEEE.numeric_std.ALL;

entity Instr_Memory is
  GENERIC (N:     NATURAL:= 32);  -- Width of inputs.
  port (address : in std_logic_vector(N-1 downto 0);			
		data    : out std_logic_vector(N-1 downto 0));
end Instr_Memory;

architecture behavioral of Instr_Memory is
signal addr : integer range 0 to 4*50760;  
 
begin
addr <= to_integer(unsigned(address));
   process(addr) 
	begin
      case addr is 
       when 4*0    => data <= "10000100001000000000000000000001"; -- addi r01,r00,1
       when 4*1    => data <= "00000000000000000000000000000000"; -- nop
       when 4*2    => data <= "00000000000000000000000000000000"; -- nop
       when 4*3    => data <= "00000000000000000000000000000000"; -- nop
       when 4*4    => data <= "00000000000000000000000000000000"; -- nop
       when 4*5    => data <= "00000000000000000000000000000000"; -- nop
       when 4*6    => data <= "10000100010000010000000000000010"; -- addi r02,r01,2
       when 4*7    => data <= "00000000000000000000000000000000"; -- nop
       when 4*8    => data <= "00000000000000000000000000000000"; -- nop
       when 4*9    => data <= "00000000000000000000000000000000"; -- nop
       when 4*10   => data <= "00000000000000000000000000000000"; -- nop
       when 4*11   => data <= "00000000000000000000000000000000"; -- nop
       when 4*12   => data <= "10000100011000100000000000000011"; -- addi r03,r02,3
       when 4*13   => data <= "00000000000000000000000000000000"; -- nop
       when 4*14   => data <= "00000000000000000000000000000000"; -- nop
       when 4*15   => data <= "00000000000000000000000000000000"; -- nop
       when 4*16   => data <= "00000000000000000000000000000000"; -- nop
       when 4*17   => data <= "00000000000000000000000000000000"; -- nop
       when 4*18   => data <= "10000100100000110000000000000100"; -- addi r04,r03,4
       when 4*19   => data <= "00000000000000000000000000000000"; -- nop
       when 4*20   => data <= "00000000000000000000000000000000"; -- nop
       when 4*21   => data <= "00000000000000000000000000000000"; -- nop
       when 4*22   => data <= "00000000000000000000000000000000"; -- nop
       when 4*23   => data <= "00000000000000000000000000000000"; -- nop
       when 4*24   => data <= "00000011111000010001100000100000"; -- add r31,r01,r03
       when 4*25   => data <= "00000000000000000000000000000000"; -- nop
       when 4*26   => data <= "00000000000000000000000000000000"; -- nop
       when 4*27   => data <= "00000000000000000000000000000000"; -- nop
       when 4*28   => data <= "00000000000000000000000000000000"; -- nop
       when 4*29   => data <= "00000000000000000000000000000000"; -- nop
       when 4*30   => data <= "00000011110111110000100000100000"; -- add r30,r31,r01
       when 4*31   => data <= "00000000000000000000000000000000"; -- nop
       when 4*32   => data <= "00000000000000000000000000000000"; -- nop
       when 4*33   => data <= "00000000000000000000000000000000"; -- nop
       when 4*34   => data <= "00000000000000000000000000000000"; -- nop
       when 4*35   => data <= "00000000000000000000000000000000"; -- nop
       when 4*36   => data <= "00000011111111110001000000100010"; -- sub r31,r31,r02
       when 4*37   => data <= "00000000000000000000000000000000"; -- nop
       when 4*38   => data <= "00000000000000000000000000000000"; -- nop
       when 4*39   => data <= "00000000000000000000000000000000"; -- nop
       when 4*40   => data <= "00000000000000000000000000000000"; -- nop
       when 4*41   => data <= "00000000000000000000000000000000"; -- nop
       when 4*42   => data <= "11000000001000000000000000000001"; -- sb r01,r00,1
       when 4*43   => data <= "11000000010000000000000000000010"; -- sb r02,r00,2
       when 4*44   => data <= "00000000000000000000000000000000"; -- nop
       when 4*45   => data <= "00000000000000000000000000000000"; -- nop
       when 4*46   => data <= "00000000000000000000000000000000"; -- nop
       when 4*47   => data <= "00000000000000000000000000000000"; -- nop
       when 4*48   => data <= "00000000000000000000000000000000"; -- nop
       when 4*49   => data <= "00000000000000000000000000000000"; -- nop
       when 4*50   => data <= "00000000000000000000000000000000"; -- nop
       when 4*51   => data <= "00000000000000000000000000000000"; -- nop
       when 4*52   => data <= "00000000000000000000000000000000"; -- nop
       when 4*53   => data <= "00000000000000000000000000000000"; -- nop
       when 4*54   => data <= "10000100001000000000000000000001"; -- addi r01,r00,1
       when 4*55   => data <= "10000100010000000000000000000010"; -- addi r02,r00,2
       when 4*56   => data <= "10000100011000000000000000000011"; -- addi r03,r00,3
       when 4*57   => data <= "10000100100000000000000000000100"; -- addi r04,r00,4
       when 4*58   => data <= "00000000000000000000000000000000"; -- nop
       when 4*59   => data <= "00000000000000000000000000000000"; -- nop
       when 4*60   => data <= "00000000000000000000000000000000"; -- nop
       when 4*61   => data <= "00000000000000000000000000000000"; -- nop
       when 4*62   => data <= "00000000000000000000000000000000"; -- nop
       when 4*63   => data <= "00000011111000100001000000100100"; -- mult r31,r02,r02
       when 4*64   => data <= "00000000000000000000000000000000"; -- nop
       when 4*65   => data <= "00000000000000000000000000000000"; -- nop
       when 4*66   => data <= "00000000000000000000000000000000"; -- nop
       when 4*67   => data <= "00000000000000000000000000000000"; -- nop
       when 4*68   => data <= "00000000000000000000000000000000"; -- nop
       when 4*69   => data <= "00000011111000100001100000100100"; -- mult r31,r02,r03
       when 4*70   => data <= "00000000000000000000000000000000"; -- nop
       when 4*71   => data <= "00000000000000000000000000000000"; -- nop
       when 4*72   => data <= "00000000000000000000000000000000"; -- nop
       when 4*73   => data <= "00000000000000000000000000000000"; -- nop
       when 4*74   => data <= "00000000000000000000000000000000"; -- nop
       when 4*75   => data <= "10000000001000000000000000000001"; -- lb r01,r00,1
       when 4*76   => data <= "10000000010000000000000000000010"; -- lb r02,r00,2
	    when others => data <= "00000000000000000000000000000000"; 
       end case;
	end process;
end behavioral;
