library ieee;
use ieee.std_logic_1164.all;
USE IEEE.numeric_std.ALL;

entity Instr_Memory is
  GENERIC (N:     NATURAL:= 32);  -- Width of inputs.
  port (address : in std_logic_vector(N-1 downto 0);			
		data    : out std_logic_vector(N-1 downto 0));
end Instr_Memory;

architecture behavioral of Instr_Memory is
signal addr : integer range 0 to 4*50760;  
 
begin
addr <= to_integer(unsigned(address));
   process(addr) 
	begin
      case addr is 
       when 4*0    => data <= "00000000000000000000000000000000"; -- nop
       when 4*1    => data <= "00000000000000000000000000000000"; -- nop
       when 4*2    => data <= "00000000000000000000000000000000"; -- nop
       when 4*3    => data <= "00000000000000000000000000000000"; -- nop
       when 4*4    => data <= "00000000000000000000000000000000"; -- nop
       when 4*5    => data <= "11000010100000000000000000000101"; -- sb r20,r00,5
       when 4*6    => data <= "00000000000000000000000000000000"; -- nop
       when 4*7    => data <= "00000000000000000000000000000000"; -- nop
       when 4*8    => data <= "00000000000000000000000000000000"; -- nop
       when 4*9    => data <= "00000000000000000000000000000000"; -- nop
       when 4*10   => data <= "00000000000000000000000000000000"; -- nop
       when 4*11   => data <= "10000001010000000000000000000101"; -- lb r10,r00,5
       when 4*12   => data <= "00000000000000000000000000000000"; -- nop
       when 4*13   => data <= "00000000000000000000000000000000"; -- nop
       when 4*14   => data <= "00000000000000000000000000000000"; -- nop
       when 4*15   => data <= "00000000000000000000000000000000"; -- nop
       when 4*16   => data <= "00000000000000000000000000000000"; -- nop
       when 4*17   => data <= "10000001010000000000000000000001"; -- lb r10,r00,1
       when 4*18   => data <= "00000000000000000000000000000000"; -- nop
       when 4*19   => data <= "00000000000000000000000000000000"; -- nop
       when 4*20   => data <= "00000000000000000000000000000000"; -- nop
       when 4*21   => data <= "00000000000000000000000000000000"; -- nop
       when 4*22   => data <= "00000000000000000000000000000000"; -- nop
       when 4*23   => data <= "00001001010001100000000000111010"; -- beq r10,r06,READMEM
       when 4*24   => data <= "00000000000000000000000000000000"; -- nop
       when 4*25   => data <= "00000000000000000000000000000000"; -- nop
       when 4*26   => data <= "00000000000000000000000000000000"; -- nop
       when 4*27   => data <= "00000000000000000000000000000000"; -- nop
       when 4*28   => data <= "00000000000000000000000000000000"; -- nop
       when 4*29   => data <= "00000100000000000000000000001100"; -- jmp READUART
       when 4*30   => data <= "00000000000000000000000000000000"; -- nop
       when 4*31   => data <= "00000000000000000000000000000000"; -- nop
       when 4*32   => data <= "00000000000000000000000000000000"; -- nop
       when 4*33   => data <= "00001000000010100000000000001100"; -- beq r00,r10,READUART
       when 4*34   => data <= "00000000000000000000000000000000"; -- nop
       when 4*35   => data <= "00000000000000000000000000000000"; -- nop
       when 4*36   => data <= "00000000000000000000000000000000"; -- nop
       when 4*37   => data <= "00000000000000000000000000000000"; -- nop
       when 4*38   => data <= "00000000000000000000000000000000"; -- nop
       when 4*39   => data <= "11000001010000010000000000000010"; -- sb r10,r01,2
       when 4*40   => data <= "00001000001001010000000000111010"; -- beq r01,r05,READMEM
       when 4*41   => data <= "00000000000000000000000000000000"; -- nop
       when 4*42   => data <= "00000000000000000000000000000000"; -- nop
       when 4*43   => data <= "00000000000000000000000000000000"; -- nop
       when 4*44   => data <= "00000000000000000000000000000000"; -- nop
       when 4*45   => data <= "00000000000000000000000000000000"; -- nop
       when 4*46   => data <= "10000100001000010000000000000001"; -- addi r01,r01,1
       when 4*47   => data <= "00000000000000000000000000000000"; -- nop
       when 4*48   => data <= "00000000000000000000000000000000"; -- nop
       when 4*49   => data <= "00000000000000000000000000000000"; -- nop
       when 4*50   => data <= "00000000000000000000000000000000"; -- nop
       when 4*51   => data <= "00000000000000000000000000000000"; -- nop
       when 4*52   => data <= "00000100000000000000000000001100"; -- jmp READUART
       when 4*53   => data <= "00000000000000000000000000000000"; -- nop
       when 4*54   => data <= "00000000000000000000000000000000"; -- nop
       when 4*55   => data <= "00000000000000000000000000000000"; -- nop
       when 4*56   => data <= "00000000000000000000000000000000"; -- nop
       when 4*57   => data <= "00000000000000000000000000000000"; -- nop
       when 4*58   => data <= "00000000000000000000000000000000"; -- nop
       when 4*59   => data <= "00000000000000000000000000000000"; -- nop
       when 4*60   => data <= "00000000000000000000000000000000"; -- nop
       when 4*61   => data <= "00000000000000000000000000000000"; -- nop
       when 4*62   => data <= "00000000000000000000000000000000"; -- nop
       when 4*63   => data <= "10000001011000010000000000000010"; -- lb r11,r01,2
       when 4*64   => data <= "00000000000000000000000000000000"; -- nop
       when 4*65   => data <= "00000000000000000000000000000000"; -- nop
       when 4*66   => data <= "00000000000000000000000000000000"; -- nop
       when 4*67   => data <= "00000000000000000000000000000000"; -- nop
       when 4*68   => data <= "00000000000000000000000000000000"; -- nop
       when 4*69   => data <= "11000001011000000000000000000000"; -- sb r11,r00,0
       when 4*70   => data <= "00000000000000000000000000000000"; -- nop
       when 4*71   => data <= "00000000000000000000000000000000"; -- nop
       when 4*72   => data <= "00000000000000000000000000000000"; -- nop
       when 4*73   => data <= "00000000000000000000000000000000"; -- nop
       when 4*74   => data <= "00000000000000000000000000000000"; -- nop
       when 4*75   => data <= "00000100000000000000000001000000"; -- jmp OUTPUT
       when 4*76   => data <= "00000000000000000000000000000000"; -- nop
       when 4*77   => data <= "00000000000000000000000000000000"; -- nop
       when 4*78   => data <= "00000000000000000000000000000000"; -- nop
       when 4*79   => data <= "00000000000000000000000000000000"; -- nop
       when 4*80   => data <= "00000000000000000000000000000000"; -- nop
       when 4*81   => data <= "00001000001000000000000001011110"; -- beq r01,r00,END
       when 4*82   => data <= "00000000000000000000000000000000"; -- nop
       when 4*83   => data <= "00000000000000000000000000000000"; -- nop
       when 4*84   => data <= "00000000000000000000000000000000"; -- nop
       when 4*85   => data <= "00000000000000000000000000000000"; -- nop
       when 4*86   => data <= "00000000000000000000000000000000"; -- nop
       when 4*87   => data <= "00000000001000010010000000100010"; -- sub r01,r01,r04
       when 4*88   => data <= "00000000000000000000000000000000"; -- nop
       when 4*89   => data <= "00000000000000000000000000000000"; -- nop
       when 4*90   => data <= "00000000000000000000000000000000"; -- nop
       when 4*91   => data <= "00000000000000000000000000000000"; -- nop
       when 4*92   => data <= "00000000000000000000000000000000"; -- nop
       when 4*93   => data <= "00000100000000000000000000111010"; -- jmp READMEM
       when 4*94   => data <= "00000000000000000000000000000000"; -- nop
       when 4*95   => data <= "00000000000000000000000000000000"; -- nop
       when 4*96   => data <= "00000000000000000000000000000000"; -- nop
       when 4*97   => data <= "00000000000000000000000000000000"; -- nop
       when 4*98   => data <= "00000000000000000000000000000000"; -- nop
	    when others => data <= "00000000000000000000000000000000"; 
       end case;
	end process;
end behavioral;
